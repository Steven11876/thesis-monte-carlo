
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_SABR.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_SABR.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_SABR.ap_done;
    assign module_intf_1.ap_continue = AESL_inst_SABR.ap_continue;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_ready;
    assign module_intf_49.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_done;
    assign module_intf_49.ap_continue = 1'b1;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_start;
    assign module_intf_50.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_ready;
    assign module_intf_50.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_done;
    assign module_intf_50.ap_continue = 1'b1;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_start;
    assign module_intf_53.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_ready;
    assign module_intf_53.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_done;
    assign module_intf_53.ap_continue = 1'b1;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_start;
    assign module_intf_54.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_ready;
    assign module_intf_54.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_done;
    assign module_intf_54.ap_continue = 1'b1;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_start;
    assign module_intf_55.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_ready;
    assign module_intf_55.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_done;
    assign module_intf_55.ap_continue = 1'b1;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_start;
    assign module_intf_56.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_ready;
    assign module_intf_56.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_done;
    assign module_intf_56.ap_continue = 1'b1;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_start;
    assign module_intf_57.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_ready;
    assign module_intf_57.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_done;
    assign module_intf_57.ap_continue = 1'b1;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_start;
    assign module_intf_58.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_ready;
    assign module_intf_58.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_done;
    assign module_intf_58.ap_continue = 1'b1;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_start;
    assign module_intf_59.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_ready;
    assign module_intf_59.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_done;
    assign module_intf_59.ap_continue = 1'b1;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_start;
    assign module_intf_60.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_ready;
    assign module_intf_60.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_done;
    assign module_intf_60.ap_continue = 1'b1;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_start;
    assign module_intf_61.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_ready;
    assign module_intf_61.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_done;
    assign module_intf_61.ap_continue = 1'b1;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_start;
    assign module_intf_62.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_ready;
    assign module_intf_62.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_done;
    assign module_intf_62.ap_continue = 1'b1;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_start;
    assign module_intf_63.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_ready;
    assign module_intf_63.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_done;
    assign module_intf_63.ap_continue = 1'b1;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_start;
    assign module_intf_64.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_ready;
    assign module_intf_64.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_done;
    assign module_intf_64.ap_continue = 1'b1;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_start;
    assign module_intf_65.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_ready;
    assign module_intf_65.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_done;
    assign module_intf_65.ap_continue = 1'b1;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_start;
    assign module_intf_66.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_ready;
    assign module_intf_66.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_done;
    assign module_intf_66.ap_continue = 1'b1;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_start;
    assign module_intf_67.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_ready;
    assign module_intf_67.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_done;
    assign module_intf_67.ap_continue = 1'b1;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;
    nodf_module_intf module_intf_68(clock,reset);
    assign module_intf_68.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_start;
    assign module_intf_68.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_ready;
    assign module_intf_68.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_done;
    assign module_intf_68.ap_continue = 1'b1;
    assign module_intf_68.finish = finish;
    csv_file_dump mstatus_csv_dumper_68;
    nodf_module_monitor module_monitor_68;
    nodf_module_intf module_intf_69(clock,reset);
    assign module_intf_69.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_start;
    assign module_intf_69.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_ready;
    assign module_intf_69.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_done;
    assign module_intf_69.ap_continue = 1'b1;
    assign module_intf_69.finish = finish;
    csv_file_dump mstatus_csv_dumper_69;
    nodf_module_monitor module_monitor_69;
    nodf_module_intf module_intf_70(clock,reset);
    assign module_intf_70.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_start;
    assign module_intf_70.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_ready;
    assign module_intf_70.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_done;
    assign module_intf_70.ap_continue = 1'b1;
    assign module_intf_70.finish = finish;
    csv_file_dump mstatus_csv_dumper_70;
    nodf_module_monitor module_monitor_70;
    nodf_module_intf module_intf_71(clock,reset);
    assign module_intf_71.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_start;
    assign module_intf_71.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_ready;
    assign module_intf_71.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_done;
    assign module_intf_71.ap_continue = 1'b1;
    assign module_intf_71.finish = finish;
    csv_file_dump mstatus_csv_dumper_71;
    nodf_module_monitor module_monitor_71;
    nodf_module_intf module_intf_72(clock,reset);
    assign module_intf_72.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_start;
    assign module_intf_72.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_ready;
    assign module_intf_72.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_done;
    assign module_intf_72.ap_continue = 1'b1;
    assign module_intf_72.finish = finish;
    csv_file_dump mstatus_csv_dumper_72;
    nodf_module_monitor module_monitor_72;
    nodf_module_intf module_intf_73(clock,reset);
    assign module_intf_73.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_start;
    assign module_intf_73.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_ready;
    assign module_intf_73.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_done;
    assign module_intf_73.ap_continue = 1'b1;
    assign module_intf_73.finish = finish;
    csv_file_dump mstatus_csv_dumper_73;
    nodf_module_monitor module_monitor_73;
    nodf_module_intf module_intf_74(clock,reset);
    assign module_intf_74.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_start;
    assign module_intf_74.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_ready;
    assign module_intf_74.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_done;
    assign module_intf_74.ap_continue = 1'b1;
    assign module_intf_74.finish = finish;
    csv_file_dump mstatus_csv_dumper_74;
    nodf_module_monitor module_monitor_74;
    nodf_module_intf module_intf_75(clock,reset);
    assign module_intf_75.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_start;
    assign module_intf_75.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_ready;
    assign module_intf_75.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_done;
    assign module_intf_75.ap_continue = 1'b1;
    assign module_intf_75.finish = finish;
    csv_file_dump mstatus_csv_dumper_75;
    nodf_module_monitor module_monitor_75;
    nodf_module_intf module_intf_76(clock,reset);
    assign module_intf_76.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_start;
    assign module_intf_76.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_ready;
    assign module_intf_76.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_done;
    assign module_intf_76.ap_continue = 1'b1;
    assign module_intf_76.finish = finish;
    csv_file_dump mstatus_csv_dumper_76;
    nodf_module_monitor module_monitor_76;
    nodf_module_intf module_intf_77(clock,reset);
    assign module_intf_77.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_start;
    assign module_intf_77.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_ready;
    assign module_intf_77.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_done;
    assign module_intf_77.ap_continue = 1'b1;
    assign module_intf_77.finish = finish;
    csv_file_dump mstatus_csv_dumper_77;
    nodf_module_monitor module_monitor_77;
    nodf_module_intf module_intf_78(clock,reset);
    assign module_intf_78.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_start;
    assign module_intf_78.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_ready;
    assign module_intf_78.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_done;
    assign module_intf_78.ap_continue = 1'b1;
    assign module_intf_78.finish = finish;
    csv_file_dump mstatus_csv_dumper_78;
    nodf_module_monitor module_monitor_78;
    nodf_module_intf module_intf_79(clock,reset);
    assign module_intf_79.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_start;
    assign module_intf_79.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_ready;
    assign module_intf_79.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_done;
    assign module_intf_79.ap_continue = 1'b1;
    assign module_intf_79.finish = finish;
    csv_file_dump mstatus_csv_dumper_79;
    nodf_module_monitor module_monitor_79;
    nodf_module_intf module_intf_80(clock,reset);
    assign module_intf_80.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_start;
    assign module_intf_80.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_ready;
    assign module_intf_80.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_done;
    assign module_intf_80.ap_continue = 1'b1;
    assign module_intf_80.finish = finish;
    csv_file_dump mstatus_csv_dumper_80;
    nodf_module_monitor module_monitor_80;
    nodf_module_intf module_intf_81(clock,reset);
    assign module_intf_81.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_start;
    assign module_intf_81.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_ready;
    assign module_intf_81.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_done;
    assign module_intf_81.ap_continue = 1'b1;
    assign module_intf_81.finish = finish;
    csv_file_dump mstatus_csv_dumper_81;
    nodf_module_monitor module_monitor_81;
    nodf_module_intf module_intf_82(clock,reset);
    assign module_intf_82.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_start;
    assign module_intf_82.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_ready;
    assign module_intf_82.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_done;
    assign module_intf_82.ap_continue = 1'b1;
    assign module_intf_82.finish = finish;
    csv_file_dump mstatus_csv_dumper_82;
    nodf_module_monitor module_monitor_82;
    nodf_module_intf module_intf_83(clock,reset);
    assign module_intf_83.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_start;
    assign module_intf_83.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_ready;
    assign module_intf_83.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_done;
    assign module_intf_83.ap_continue = 1'b1;
    assign module_intf_83.finish = finish;
    csv_file_dump mstatus_csv_dumper_83;
    nodf_module_monitor module_monitor_83;
    nodf_module_intf module_intf_84(clock,reset);
    assign module_intf_84.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_start;
    assign module_intf_84.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_ready;
    assign module_intf_84.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_done;
    assign module_intf_84.ap_continue = 1'b1;
    assign module_intf_84.finish = finish;
    csv_file_dump mstatus_csv_dumper_84;
    nodf_module_monitor module_monitor_84;
    nodf_module_intf module_intf_85(clock,reset);
    assign module_intf_85.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_start;
    assign module_intf_85.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_ready;
    assign module_intf_85.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_done;
    assign module_intf_85.ap_continue = 1'b1;
    assign module_intf_85.finish = finish;
    csv_file_dump mstatus_csv_dumper_85;
    nodf_module_monitor module_monitor_85;
    nodf_module_intf module_intf_86(clock,reset);
    assign module_intf_86.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_start;
    assign module_intf_86.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_ready;
    assign module_intf_86.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_done;
    assign module_intf_86.ap_continue = 1'b1;
    assign module_intf_86.finish = finish;
    csv_file_dump mstatus_csv_dumper_86;
    nodf_module_monitor module_monitor_86;
    nodf_module_intf module_intf_87(clock,reset);
    assign module_intf_87.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_start;
    assign module_intf_87.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_ready;
    assign module_intf_87.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_done;
    assign module_intf_87.ap_continue = 1'b1;
    assign module_intf_87.finish = finish;
    csv_file_dump mstatus_csv_dumper_87;
    nodf_module_monitor module_monitor_87;
    nodf_module_intf module_intf_88(clock,reset);
    assign module_intf_88.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_start;
    assign module_intf_88.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_ready;
    assign module_intf_88.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_done;
    assign module_intf_88.ap_continue = 1'b1;
    assign module_intf_88.finish = finish;
    csv_file_dump mstatus_csv_dumper_88;
    nodf_module_monitor module_monitor_88;
    nodf_module_intf module_intf_89(clock,reset);
    assign module_intf_89.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_start;
    assign module_intf_89.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_ready;
    assign module_intf_89.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_done;
    assign module_intf_89.ap_continue = 1'b1;
    assign module_intf_89.finish = finish;
    csv_file_dump mstatus_csv_dumper_89;
    nodf_module_monitor module_monitor_89;
    nodf_module_intf module_intf_90(clock,reset);
    assign module_intf_90.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_start;
    assign module_intf_90.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_ready;
    assign module_intf_90.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_done;
    assign module_intf_90.ap_continue = 1'b1;
    assign module_intf_90.finish = finish;
    csv_file_dump mstatus_csv_dumper_90;
    nodf_module_monitor module_monitor_90;
    nodf_module_intf module_intf_91(clock,reset);
    assign module_intf_91.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_start;
    assign module_intf_91.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_ready;
    assign module_intf_91.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_done;
    assign module_intf_91.ap_continue = 1'b1;
    assign module_intf_91.finish = finish;
    csv_file_dump mstatus_csv_dumper_91;
    nodf_module_monitor module_monitor_91;
    nodf_module_intf module_intf_92(clock,reset);
    assign module_intf_92.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_start;
    assign module_intf_92.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_ready;
    assign module_intf_92.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_done;
    assign module_intf_92.ap_continue = 1'b1;
    assign module_intf_92.finish = finish;
    csv_file_dump mstatus_csv_dumper_92;
    nodf_module_monitor module_monitor_92;
    nodf_module_intf module_intf_93(clock,reset);
    assign module_intf_93.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_start;
    assign module_intf_93.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_ready;
    assign module_intf_93.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_done;
    assign module_intf_93.ap_continue = 1'b1;
    assign module_intf_93.finish = finish;
    csv_file_dump mstatus_csv_dumper_93;
    nodf_module_monitor module_monitor_93;
    nodf_module_intf module_intf_94(clock,reset);
    assign module_intf_94.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_start;
    assign module_intf_94.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_ready;
    assign module_intf_94.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_done;
    assign module_intf_94.ap_continue = 1'b1;
    assign module_intf_94.finish = finish;
    csv_file_dump mstatus_csv_dumper_94;
    nodf_module_monitor module_monitor_94;
    nodf_module_intf module_intf_95(clock,reset);
    assign module_intf_95.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_start;
    assign module_intf_95.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_ready;
    assign module_intf_95.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_done;
    assign module_intf_95.ap_continue = 1'b1;
    assign module_intf_95.finish = finish;
    csv_file_dump mstatus_csv_dumper_95;
    nodf_module_monitor module_monitor_95;
    nodf_module_intf module_intf_96(clock,reset);
    assign module_intf_96.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_start;
    assign module_intf_96.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_ready;
    assign module_intf_96.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_done;
    assign module_intf_96.ap_continue = 1'b1;
    assign module_intf_96.finish = finish;
    csv_file_dump mstatus_csv_dumper_96;
    nodf_module_monitor module_monitor_96;
    nodf_module_intf module_intf_97(clock,reset);
    assign module_intf_97.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_start;
    assign module_intf_97.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_ready;
    assign module_intf_97.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_done;
    assign module_intf_97.ap_continue = 1'b1;
    assign module_intf_97.finish = finish;
    csv_file_dump mstatus_csv_dumper_97;
    nodf_module_monitor module_monitor_97;
    nodf_module_intf module_intf_98(clock,reset);
    assign module_intf_98.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_start;
    assign module_intf_98.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_ready;
    assign module_intf_98.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_done;
    assign module_intf_98.ap_continue = 1'b1;
    assign module_intf_98.finish = finish;
    csv_file_dump mstatus_csv_dumper_98;
    nodf_module_monitor module_monitor_98;
    nodf_module_intf module_intf_99(clock,reset);
    assign module_intf_99.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_start;
    assign module_intf_99.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_ready;
    assign module_intf_99.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_done;
    assign module_intf_99.ap_continue = 1'b1;
    assign module_intf_99.finish = finish;
    csv_file_dump mstatus_csv_dumper_99;
    nodf_module_monitor module_monitor_99;
    nodf_module_intf module_intf_100(clock,reset);
    assign module_intf_100.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_start;
    assign module_intf_100.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_ready;
    assign module_intf_100.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_done;
    assign module_intf_100.ap_continue = 1'b1;
    assign module_intf_100.finish = finish;
    csv_file_dump mstatus_csv_dumper_100;
    nodf_module_monitor module_monitor_100;
    nodf_module_intf module_intf_101(clock,reset);
    assign module_intf_101.ap_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_start;
    assign module_intf_101.ap_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_ready;
    assign module_intf_101.ap_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_done;
    assign module_intf_101.ap_continue = 1'b1;
    assign module_intf_101.finish = finish;
    csv_file_dump mstatus_csv_dumper_101;
    nodf_module_monitor module_monitor_101;
    nodf_module_intf module_intf_102(clock,reset);
    assign module_intf_102.ap_start = AESL_inst_SABR.grp_pow_generic_double_s_fu_28633.ap_start;
    assign module_intf_102.ap_ready = AESL_inst_SABR.grp_pow_generic_double_s_fu_28633.ap_ready;
    assign module_intf_102.ap_done = AESL_inst_SABR.grp_pow_generic_double_s_fu_28633.ap_done;
    assign module_intf_102.ap_continue = 1'b1;
    assign module_intf_102.finish = finish;
    csv_file_dump mstatus_csv_dumper_102;
    nodf_module_monitor module_monitor_102;

    upc_loop_intf#(34) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_1.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_3_fu_10070.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(34) upc_loop_monitor_1;
    upc_loop_intf#(34) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_2.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_31_fu_10113.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(34) upc_loop_monitor_2;
    upc_loop_intf#(34) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_3.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_32_fu_10155.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(34) upc_loop_monitor_3;
    upc_loop_intf#(34) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_4.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_33_fu_10197.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(34) upc_loop_monitor_4;
    upc_loop_intf#(34) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_5.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_34_fu_10239.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(34) upc_loop_monitor_5;
    upc_loop_intf#(34) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_6.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_35_fu_10281.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(34) upc_loop_monitor_6;
    upc_loop_intf#(34) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_7.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_36_fu_10323.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(34) upc_loop_monitor_7;
    upc_loop_intf#(34) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_8.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_37_fu_10365.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(34) upc_loop_monitor_8;
    upc_loop_intf#(34) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_9.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_38_fu_10407.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(34) upc_loop_monitor_9;
    upc_loop_intf#(34) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_10.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_39_fu_10449.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(34) upc_loop_monitor_10;
    upc_loop_intf#(34) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_11.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_310_fu_10491.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(34) upc_loop_monitor_11;
    upc_loop_intf#(34) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_12.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_311_fu_10533.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(34) upc_loop_monitor_12;
    upc_loop_intf#(34) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_13.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_312_fu_10575.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(34) upc_loop_monitor_13;
    upc_loop_intf#(34) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_14.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_313_fu_10617.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(34) upc_loop_monitor_14;
    upc_loop_intf#(34) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_15.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_314_fu_10659.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(34) upc_loop_monitor_15;
    upc_loop_intf#(34) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_16.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_315_fu_10701.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(34) upc_loop_monitor_16;
    upc_loop_intf#(34) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_17.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_316_fu_10743.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b1;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(34) upc_loop_monitor_17;
    upc_loop_intf#(34) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_18.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_18.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_18.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_317_fu_10785.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b1;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(34) upc_loop_monitor_18;
    upc_loop_intf#(34) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_19.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_318_fu_10827.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b1;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(34) upc_loop_monitor_19;
    upc_loop_intf#(34) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_20.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_319_fu_10869.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b1;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(34) upc_loop_monitor_20;
    upc_loop_intf#(34) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_21.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_320_fu_10911.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b1;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(34) upc_loop_monitor_21;
    upc_loop_intf#(34) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_22.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_22.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_22.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_321_fu_10953.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b1;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(34) upc_loop_monitor_22;
    upc_loop_intf#(34) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_23.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_322_fu_10995.ap_done_int;
    assign upc_loop_intf_23.loop_continue = 1'b1;
    assign upc_loop_intf_23.quit_at_end = 1'b1;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(34) upc_loop_monitor_23;
    upc_loop_intf#(34) upc_loop_intf_24(clock,reset);
    assign upc_loop_intf_24.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_CS_fsm;
    assign upc_loop_intf_24.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_24.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_24.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_24.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_24.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_24.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_24.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_start;
    assign upc_loop_intf_24.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_ready;
    assign upc_loop_intf_24.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_323_fu_11037.ap_done_int;
    assign upc_loop_intf_24.loop_continue = 1'b1;
    assign upc_loop_intf_24.quit_at_end = 1'b1;
    assign upc_loop_intf_24.finish = finish;
    csv_file_dump upc_loop_csv_dumper_24;
    upc_loop_monitor #(34) upc_loop_monitor_24;
    upc_loop_intf#(34) upc_loop_intf_25(clock,reset);
    assign upc_loop_intf_25.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_CS_fsm;
    assign upc_loop_intf_25.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_25.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_25.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_25.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_25.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_25.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_25.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_start;
    assign upc_loop_intf_25.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_ready;
    assign upc_loop_intf_25.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_324_fu_11079.ap_done_int;
    assign upc_loop_intf_25.loop_continue = 1'b1;
    assign upc_loop_intf_25.quit_at_end = 1'b1;
    assign upc_loop_intf_25.finish = finish;
    csv_file_dump upc_loop_csv_dumper_25;
    upc_loop_monitor #(34) upc_loop_monitor_25;
    upc_loop_intf#(34) upc_loop_intf_26(clock,reset);
    assign upc_loop_intf_26.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_CS_fsm;
    assign upc_loop_intf_26.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_26.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_26.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_26.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_26.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_26.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_26.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_26.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_start;
    assign upc_loop_intf_26.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_ready;
    assign upc_loop_intf_26.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_325_fu_11121.ap_done_int;
    assign upc_loop_intf_26.loop_continue = 1'b1;
    assign upc_loop_intf_26.quit_at_end = 1'b1;
    assign upc_loop_intf_26.finish = finish;
    csv_file_dump upc_loop_csv_dumper_26;
    upc_loop_monitor #(34) upc_loop_monitor_26;
    upc_loop_intf#(34) upc_loop_intf_27(clock,reset);
    assign upc_loop_intf_27.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_CS_fsm;
    assign upc_loop_intf_27.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_27.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_27.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_27.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_27.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_start;
    assign upc_loop_intf_27.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_ready;
    assign upc_loop_intf_27.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_326_fu_11163.ap_done_int;
    assign upc_loop_intf_27.loop_continue = 1'b1;
    assign upc_loop_intf_27.quit_at_end = 1'b1;
    assign upc_loop_intf_27.finish = finish;
    csv_file_dump upc_loop_csv_dumper_27;
    upc_loop_monitor #(34) upc_loop_monitor_27;
    upc_loop_intf#(34) upc_loop_intf_28(clock,reset);
    assign upc_loop_intf_28.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_CS_fsm;
    assign upc_loop_intf_28.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_28.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_28.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_28.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_28.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_28.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_28.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_28.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_start;
    assign upc_loop_intf_28.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_ready;
    assign upc_loop_intf_28.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_327_fu_11205.ap_done_int;
    assign upc_loop_intf_28.loop_continue = 1'b1;
    assign upc_loop_intf_28.quit_at_end = 1'b1;
    assign upc_loop_intf_28.finish = finish;
    csv_file_dump upc_loop_csv_dumper_28;
    upc_loop_monitor #(34) upc_loop_monitor_28;
    upc_loop_intf#(34) upc_loop_intf_29(clock,reset);
    assign upc_loop_intf_29.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_CS_fsm;
    assign upc_loop_intf_29.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_29.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_29.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_29.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_29.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_29.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_start;
    assign upc_loop_intf_29.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_ready;
    assign upc_loop_intf_29.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_328_fu_11247.ap_done_int;
    assign upc_loop_intf_29.loop_continue = 1'b1;
    assign upc_loop_intf_29.quit_at_end = 1'b1;
    assign upc_loop_intf_29.finish = finish;
    csv_file_dump upc_loop_csv_dumper_29;
    upc_loop_monitor #(34) upc_loop_monitor_29;
    upc_loop_intf#(34) upc_loop_intf_30(clock,reset);
    assign upc_loop_intf_30.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_CS_fsm;
    assign upc_loop_intf_30.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_30.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_30.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_30.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_30.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_30.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_30.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_30.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_start;
    assign upc_loop_intf_30.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_ready;
    assign upc_loop_intf_30.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_329_fu_11289.ap_done_int;
    assign upc_loop_intf_30.loop_continue = 1'b1;
    assign upc_loop_intf_30.quit_at_end = 1'b1;
    assign upc_loop_intf_30.finish = finish;
    csv_file_dump upc_loop_csv_dumper_30;
    upc_loop_monitor #(34) upc_loop_monitor_30;
    upc_loop_intf#(34) upc_loop_intf_31(clock,reset);
    assign upc_loop_intf_31.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_CS_fsm;
    assign upc_loop_intf_31.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_31.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_31.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_31.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_31.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_31.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_31.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_start;
    assign upc_loop_intf_31.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_ready;
    assign upc_loop_intf_31.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_330_fu_11331.ap_done_int;
    assign upc_loop_intf_31.loop_continue = 1'b1;
    assign upc_loop_intf_31.quit_at_end = 1'b1;
    assign upc_loop_intf_31.finish = finish;
    csv_file_dump upc_loop_csv_dumper_31;
    upc_loop_monitor #(34) upc_loop_monitor_31;
    upc_loop_intf#(34) upc_loop_intf_32(clock,reset);
    assign upc_loop_intf_32.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_CS_fsm;
    assign upc_loop_intf_32.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_32.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_32.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_32.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_32.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_32.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_32.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_32.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_start;
    assign upc_loop_intf_32.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_ready;
    assign upc_loop_intf_32.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_331_fu_11373.ap_done_int;
    assign upc_loop_intf_32.loop_continue = 1'b1;
    assign upc_loop_intf_32.quit_at_end = 1'b1;
    assign upc_loop_intf_32.finish = finish;
    csv_file_dump upc_loop_csv_dumper_32;
    upc_loop_monitor #(34) upc_loop_monitor_32;
    upc_loop_intf#(34) upc_loop_intf_33(clock,reset);
    assign upc_loop_intf_33.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_CS_fsm;
    assign upc_loop_intf_33.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_33.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_33.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_33.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_33.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_33.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_start;
    assign upc_loop_intf_33.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_ready;
    assign upc_loop_intf_33.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_332_fu_11415.ap_done_int;
    assign upc_loop_intf_33.loop_continue = 1'b1;
    assign upc_loop_intf_33.quit_at_end = 1'b1;
    assign upc_loop_intf_33.finish = finish;
    csv_file_dump upc_loop_csv_dumper_33;
    upc_loop_monitor #(34) upc_loop_monitor_33;
    upc_loop_intf#(34) upc_loop_intf_34(clock,reset);
    assign upc_loop_intf_34.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_CS_fsm;
    assign upc_loop_intf_34.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_34.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_34.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_34.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_34.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_34.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_start;
    assign upc_loop_intf_34.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_ready;
    assign upc_loop_intf_34.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_333_fu_11457.ap_done_int;
    assign upc_loop_intf_34.loop_continue = 1'b1;
    assign upc_loop_intf_34.quit_at_end = 1'b1;
    assign upc_loop_intf_34.finish = finish;
    csv_file_dump upc_loop_csv_dumper_34;
    upc_loop_monitor #(34) upc_loop_monitor_34;
    upc_loop_intf#(34) upc_loop_intf_35(clock,reset);
    assign upc_loop_intf_35.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_CS_fsm;
    assign upc_loop_intf_35.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_35.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_35.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_35.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_35.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_35.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_start;
    assign upc_loop_intf_35.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_ready;
    assign upc_loop_intf_35.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_334_fu_11499.ap_done_int;
    assign upc_loop_intf_35.loop_continue = 1'b1;
    assign upc_loop_intf_35.quit_at_end = 1'b1;
    assign upc_loop_intf_35.finish = finish;
    csv_file_dump upc_loop_csv_dumper_35;
    upc_loop_monitor #(34) upc_loop_monitor_35;
    upc_loop_intf#(34) upc_loop_intf_36(clock,reset);
    assign upc_loop_intf_36.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_CS_fsm;
    assign upc_loop_intf_36.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_36.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_36.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_36.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_36.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_36.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_start;
    assign upc_loop_intf_36.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_ready;
    assign upc_loop_intf_36.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_335_fu_11541.ap_done_int;
    assign upc_loop_intf_36.loop_continue = 1'b1;
    assign upc_loop_intf_36.quit_at_end = 1'b1;
    assign upc_loop_intf_36.finish = finish;
    csv_file_dump upc_loop_csv_dumper_36;
    upc_loop_monitor #(34) upc_loop_monitor_36;
    upc_loop_intf#(34) upc_loop_intf_37(clock,reset);
    assign upc_loop_intf_37.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_CS_fsm;
    assign upc_loop_intf_37.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_37.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_37.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_37.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_37.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_37.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_37.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_37.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_start;
    assign upc_loop_intf_37.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_ready;
    assign upc_loop_intf_37.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_336_fu_11583.ap_done_int;
    assign upc_loop_intf_37.loop_continue = 1'b1;
    assign upc_loop_intf_37.quit_at_end = 1'b1;
    assign upc_loop_intf_37.finish = finish;
    csv_file_dump upc_loop_csv_dumper_37;
    upc_loop_monitor #(34) upc_loop_monitor_37;
    upc_loop_intf#(34) upc_loop_intf_38(clock,reset);
    assign upc_loop_intf_38.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_CS_fsm;
    assign upc_loop_intf_38.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_38.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_38.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_38.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_38.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_38.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_38.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_38.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_start;
    assign upc_loop_intf_38.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_ready;
    assign upc_loop_intf_38.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_337_fu_11625.ap_done_int;
    assign upc_loop_intf_38.loop_continue = 1'b1;
    assign upc_loop_intf_38.quit_at_end = 1'b1;
    assign upc_loop_intf_38.finish = finish;
    csv_file_dump upc_loop_csv_dumper_38;
    upc_loop_monitor #(34) upc_loop_monitor_38;
    upc_loop_intf#(34) upc_loop_intf_39(clock,reset);
    assign upc_loop_intf_39.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_CS_fsm;
    assign upc_loop_intf_39.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_39.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_39.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_39.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_39.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_39.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_39.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_39.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_39.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_39.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_start;
    assign upc_loop_intf_39.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_ready;
    assign upc_loop_intf_39.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_338_fu_11667.ap_done_int;
    assign upc_loop_intf_39.loop_continue = 1'b1;
    assign upc_loop_intf_39.quit_at_end = 1'b1;
    assign upc_loop_intf_39.finish = finish;
    csv_file_dump upc_loop_csv_dumper_39;
    upc_loop_monitor #(34) upc_loop_monitor_39;
    upc_loop_intf#(34) upc_loop_intf_40(clock,reset);
    assign upc_loop_intf_40.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_CS_fsm;
    assign upc_loop_intf_40.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_40.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_40.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_40.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_40.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_40.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_40.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_40.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_40.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_40.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_start;
    assign upc_loop_intf_40.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_ready;
    assign upc_loop_intf_40.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_339_fu_11709.ap_done_int;
    assign upc_loop_intf_40.loop_continue = 1'b1;
    assign upc_loop_intf_40.quit_at_end = 1'b1;
    assign upc_loop_intf_40.finish = finish;
    csv_file_dump upc_loop_csv_dumper_40;
    upc_loop_monitor #(34) upc_loop_monitor_40;
    upc_loop_intf#(34) upc_loop_intf_41(clock,reset);
    assign upc_loop_intf_41.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_CS_fsm;
    assign upc_loop_intf_41.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_41.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_41.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_41.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_41.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_41.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_41.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_41.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_41.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_41.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_start;
    assign upc_loop_intf_41.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_ready;
    assign upc_loop_intf_41.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_340_fu_11751.ap_done_int;
    assign upc_loop_intf_41.loop_continue = 1'b1;
    assign upc_loop_intf_41.quit_at_end = 1'b1;
    assign upc_loop_intf_41.finish = finish;
    csv_file_dump upc_loop_csv_dumper_41;
    upc_loop_monitor #(34) upc_loop_monitor_41;
    upc_loop_intf#(34) upc_loop_intf_42(clock,reset);
    assign upc_loop_intf_42.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_CS_fsm;
    assign upc_loop_intf_42.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_42.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_42.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_42.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_42.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_42.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_42.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_42.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_42.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_42.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_start;
    assign upc_loop_intf_42.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_ready;
    assign upc_loop_intf_42.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_341_fu_11793.ap_done_int;
    assign upc_loop_intf_42.loop_continue = 1'b1;
    assign upc_loop_intf_42.quit_at_end = 1'b1;
    assign upc_loop_intf_42.finish = finish;
    csv_file_dump upc_loop_csv_dumper_42;
    upc_loop_monitor #(34) upc_loop_monitor_42;
    upc_loop_intf#(34) upc_loop_intf_43(clock,reset);
    assign upc_loop_intf_43.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_CS_fsm;
    assign upc_loop_intf_43.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_43.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_43.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_43.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_43.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_43.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_43.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_43.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_43.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_43.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_start;
    assign upc_loop_intf_43.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_ready;
    assign upc_loop_intf_43.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_342_fu_11835.ap_done_int;
    assign upc_loop_intf_43.loop_continue = 1'b1;
    assign upc_loop_intf_43.quit_at_end = 1'b1;
    assign upc_loop_intf_43.finish = finish;
    csv_file_dump upc_loop_csv_dumper_43;
    upc_loop_monitor #(34) upc_loop_monitor_43;
    upc_loop_intf#(34) upc_loop_intf_44(clock,reset);
    assign upc_loop_intf_44.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_CS_fsm;
    assign upc_loop_intf_44.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_44.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_44.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_44.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_44.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_44.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_44.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_44.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_44.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_44.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_start;
    assign upc_loop_intf_44.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_ready;
    assign upc_loop_intf_44.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_343_fu_11877.ap_done_int;
    assign upc_loop_intf_44.loop_continue = 1'b1;
    assign upc_loop_intf_44.quit_at_end = 1'b1;
    assign upc_loop_intf_44.finish = finish;
    csv_file_dump upc_loop_csv_dumper_44;
    upc_loop_monitor #(34) upc_loop_monitor_44;
    upc_loop_intf#(34) upc_loop_intf_45(clock,reset);
    assign upc_loop_intf_45.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_CS_fsm;
    assign upc_loop_intf_45.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_45.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_45.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_45.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_45.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_45.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_45.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_45.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_45.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_45.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_start;
    assign upc_loop_intf_45.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_ready;
    assign upc_loop_intf_45.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_344_fu_11919.ap_done_int;
    assign upc_loop_intf_45.loop_continue = 1'b1;
    assign upc_loop_intf_45.quit_at_end = 1'b1;
    assign upc_loop_intf_45.finish = finish;
    csv_file_dump upc_loop_csv_dumper_45;
    upc_loop_monitor #(34) upc_loop_monitor_45;
    upc_loop_intf#(34) upc_loop_intf_46(clock,reset);
    assign upc_loop_intf_46.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_CS_fsm;
    assign upc_loop_intf_46.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_46.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_46.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_46.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_46.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_46.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_46.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_46.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_46.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_46.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_start;
    assign upc_loop_intf_46.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_ready;
    assign upc_loop_intf_46.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_345_fu_11961.ap_done_int;
    assign upc_loop_intf_46.loop_continue = 1'b1;
    assign upc_loop_intf_46.quit_at_end = 1'b1;
    assign upc_loop_intf_46.finish = finish;
    csv_file_dump upc_loop_csv_dumper_46;
    upc_loop_monitor #(34) upc_loop_monitor_46;
    upc_loop_intf#(34) upc_loop_intf_47(clock,reset);
    assign upc_loop_intf_47.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_CS_fsm;
    assign upc_loop_intf_47.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_47.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_47.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_47.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_47.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_47.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_47.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_47.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_47.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_47.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_start;
    assign upc_loop_intf_47.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_ready;
    assign upc_loop_intf_47.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_346_fu_12003.ap_done_int;
    assign upc_loop_intf_47.loop_continue = 1'b1;
    assign upc_loop_intf_47.quit_at_end = 1'b1;
    assign upc_loop_intf_47.finish = finish;
    csv_file_dump upc_loop_csv_dumper_47;
    upc_loop_monitor #(34) upc_loop_monitor_47;
    upc_loop_intf#(34) upc_loop_intf_48(clock,reset);
    assign upc_loop_intf_48.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_CS_fsm;
    assign upc_loop_intf_48.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_48.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_48.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_48.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_48.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_48.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_48.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_48.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_48.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_48.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_start;
    assign upc_loop_intf_48.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_ready;
    assign upc_loop_intf_48.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_347_fu_12045.ap_done_int;
    assign upc_loop_intf_48.loop_continue = 1'b1;
    assign upc_loop_intf_48.quit_at_end = 1'b1;
    assign upc_loop_intf_48.finish = finish;
    csv_file_dump upc_loop_csv_dumper_48;
    upc_loop_monitor #(34) upc_loop_monitor_48;
    upc_loop_intf#(34) upc_loop_intf_49(clock,reset);
    assign upc_loop_intf_49.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_CS_fsm;
    assign upc_loop_intf_49.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_49.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_49.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_49.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_49.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_49.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_49.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_49.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_49.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_49.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_start;
    assign upc_loop_intf_49.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_ready;
    assign upc_loop_intf_49.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_348_fu_12087.ap_done_int;
    assign upc_loop_intf_49.loop_continue = 1'b1;
    assign upc_loop_intf_49.quit_at_end = 1'b1;
    assign upc_loop_intf_49.finish = finish;
    csv_file_dump upc_loop_csv_dumper_49;
    upc_loop_monitor #(34) upc_loop_monitor_49;
    upc_loop_intf#(34) upc_loop_intf_50(clock,reset);
    assign upc_loop_intf_50.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_CS_fsm;
    assign upc_loop_intf_50.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_50.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_50.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_50.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_50.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_50.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_50.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_50.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_50.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_50.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_start;
    assign upc_loop_intf_50.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_ready;
    assign upc_loop_intf_50.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_349_fu_12129.ap_done_int;
    assign upc_loop_intf_50.loop_continue = 1'b1;
    assign upc_loop_intf_50.quit_at_end = 1'b1;
    assign upc_loop_intf_50.finish = finish;
    csv_file_dump upc_loop_csv_dumper_50;
    upc_loop_monitor #(34) upc_loop_monitor_50;
    upc_loop_intf#(34) upc_loop_intf_51(clock,reset);
    assign upc_loop_intf_51.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_CS_fsm;
    assign upc_loop_intf_51.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_51.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_51.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_51.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_51.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_51.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_51.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_51.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_51.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_51.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_start;
    assign upc_loop_intf_51.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_ready;
    assign upc_loop_intf_51.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_350_fu_12171.ap_done_int;
    assign upc_loop_intf_51.loop_continue = 1'b1;
    assign upc_loop_intf_51.quit_at_end = 1'b1;
    assign upc_loop_intf_51.finish = finish;
    csv_file_dump upc_loop_csv_dumper_51;
    upc_loop_monitor #(34) upc_loop_monitor_51;
    upc_loop_intf#(34) upc_loop_intf_52(clock,reset);
    assign upc_loop_intf_52.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_CS_fsm;
    assign upc_loop_intf_52.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_52.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_52.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_52.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_52.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_52.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_52.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_52.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_52.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_52.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_start;
    assign upc_loop_intf_52.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_ready;
    assign upc_loop_intf_52.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_351_fu_12213.ap_done_int;
    assign upc_loop_intf_52.loop_continue = 1'b1;
    assign upc_loop_intf_52.quit_at_end = 1'b1;
    assign upc_loop_intf_52.finish = finish;
    csv_file_dump upc_loop_csv_dumper_52;
    upc_loop_monitor #(34) upc_loop_monitor_52;
    upc_loop_intf#(34) upc_loop_intf_53(clock,reset);
    assign upc_loop_intf_53.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_CS_fsm;
    assign upc_loop_intf_53.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_53.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_53.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_53.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_53.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_53.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_53.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_53.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_53.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_53.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_start;
    assign upc_loop_intf_53.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_ready;
    assign upc_loop_intf_53.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_352_fu_12255.ap_done_int;
    assign upc_loop_intf_53.loop_continue = 1'b1;
    assign upc_loop_intf_53.quit_at_end = 1'b1;
    assign upc_loop_intf_53.finish = finish;
    csv_file_dump upc_loop_csv_dumper_53;
    upc_loop_monitor #(34) upc_loop_monitor_53;
    upc_loop_intf#(34) upc_loop_intf_54(clock,reset);
    assign upc_loop_intf_54.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_CS_fsm;
    assign upc_loop_intf_54.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_54.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_54.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_54.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_54.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_54.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_54.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_54.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_54.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_54.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_start;
    assign upc_loop_intf_54.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_ready;
    assign upc_loop_intf_54.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_353_fu_12297.ap_done_int;
    assign upc_loop_intf_54.loop_continue = 1'b1;
    assign upc_loop_intf_54.quit_at_end = 1'b1;
    assign upc_loop_intf_54.finish = finish;
    csv_file_dump upc_loop_csv_dumper_54;
    upc_loop_monitor #(34) upc_loop_monitor_54;
    upc_loop_intf#(34) upc_loop_intf_55(clock,reset);
    assign upc_loop_intf_55.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_CS_fsm;
    assign upc_loop_intf_55.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_55.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_55.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_55.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_55.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_55.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_55.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_55.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_55.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_55.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_start;
    assign upc_loop_intf_55.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_ready;
    assign upc_loop_intf_55.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_354_fu_12339.ap_done_int;
    assign upc_loop_intf_55.loop_continue = 1'b1;
    assign upc_loop_intf_55.quit_at_end = 1'b1;
    assign upc_loop_intf_55.finish = finish;
    csv_file_dump upc_loop_csv_dumper_55;
    upc_loop_monitor #(34) upc_loop_monitor_55;
    upc_loop_intf#(34) upc_loop_intf_56(clock,reset);
    assign upc_loop_intf_56.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_CS_fsm;
    assign upc_loop_intf_56.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_56.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_56.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_56.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_56.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_56.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_56.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_56.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_56.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_56.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_start;
    assign upc_loop_intf_56.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_ready;
    assign upc_loop_intf_56.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_355_fu_12381.ap_done_int;
    assign upc_loop_intf_56.loop_continue = 1'b1;
    assign upc_loop_intf_56.quit_at_end = 1'b1;
    assign upc_loop_intf_56.finish = finish;
    csv_file_dump upc_loop_csv_dumper_56;
    upc_loop_monitor #(34) upc_loop_monitor_56;
    upc_loop_intf#(34) upc_loop_intf_57(clock,reset);
    assign upc_loop_intf_57.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_CS_fsm;
    assign upc_loop_intf_57.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_57.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_57.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_57.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_57.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_57.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_57.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_57.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_57.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_57.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_start;
    assign upc_loop_intf_57.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_ready;
    assign upc_loop_intf_57.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_356_fu_12423.ap_done_int;
    assign upc_loop_intf_57.loop_continue = 1'b1;
    assign upc_loop_intf_57.quit_at_end = 1'b1;
    assign upc_loop_intf_57.finish = finish;
    csv_file_dump upc_loop_csv_dumper_57;
    upc_loop_monitor #(34) upc_loop_monitor_57;
    upc_loop_intf#(34) upc_loop_intf_58(clock,reset);
    assign upc_loop_intf_58.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_CS_fsm;
    assign upc_loop_intf_58.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_58.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_58.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_58.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_58.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_58.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_58.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_58.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_58.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_58.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_start;
    assign upc_loop_intf_58.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_ready;
    assign upc_loop_intf_58.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_357_fu_12465.ap_done_int;
    assign upc_loop_intf_58.loop_continue = 1'b1;
    assign upc_loop_intf_58.quit_at_end = 1'b1;
    assign upc_loop_intf_58.finish = finish;
    csv_file_dump upc_loop_csv_dumper_58;
    upc_loop_monitor #(34) upc_loop_monitor_58;
    upc_loop_intf#(34) upc_loop_intf_59(clock,reset);
    assign upc_loop_intf_59.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_CS_fsm;
    assign upc_loop_intf_59.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_59.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_59.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_59.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_59.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_59.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_59.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_59.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_59.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_59.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_start;
    assign upc_loop_intf_59.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_ready;
    assign upc_loop_intf_59.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_358_fu_12507.ap_done_int;
    assign upc_loop_intf_59.loop_continue = 1'b1;
    assign upc_loop_intf_59.quit_at_end = 1'b1;
    assign upc_loop_intf_59.finish = finish;
    csv_file_dump upc_loop_csv_dumper_59;
    upc_loop_monitor #(34) upc_loop_monitor_59;
    upc_loop_intf#(34) upc_loop_intf_60(clock,reset);
    assign upc_loop_intf_60.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_CS_fsm;
    assign upc_loop_intf_60.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_60.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_60.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_60.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_60.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_60.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_60.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_60.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_60.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_60.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_start;
    assign upc_loop_intf_60.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_ready;
    assign upc_loop_intf_60.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_359_fu_12549.ap_done_int;
    assign upc_loop_intf_60.loop_continue = 1'b1;
    assign upc_loop_intf_60.quit_at_end = 1'b1;
    assign upc_loop_intf_60.finish = finish;
    csv_file_dump upc_loop_csv_dumper_60;
    upc_loop_monitor #(34) upc_loop_monitor_60;
    upc_loop_intf#(34) upc_loop_intf_61(clock,reset);
    assign upc_loop_intf_61.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_CS_fsm;
    assign upc_loop_intf_61.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_61.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_61.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_61.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_61.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_61.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_61.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_61.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_61.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_61.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_start;
    assign upc_loop_intf_61.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_ready;
    assign upc_loop_intf_61.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_360_fu_12591.ap_done_int;
    assign upc_loop_intf_61.loop_continue = 1'b1;
    assign upc_loop_intf_61.quit_at_end = 1'b1;
    assign upc_loop_intf_61.finish = finish;
    csv_file_dump upc_loop_csv_dumper_61;
    upc_loop_monitor #(34) upc_loop_monitor_61;
    upc_loop_intf#(34) upc_loop_intf_62(clock,reset);
    assign upc_loop_intf_62.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_CS_fsm;
    assign upc_loop_intf_62.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_62.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_62.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_62.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_62.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_62.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_62.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_62.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_62.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_62.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_start;
    assign upc_loop_intf_62.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_ready;
    assign upc_loop_intf_62.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_361_fu_12633.ap_done_int;
    assign upc_loop_intf_62.loop_continue = 1'b1;
    assign upc_loop_intf_62.quit_at_end = 1'b1;
    assign upc_loop_intf_62.finish = finish;
    csv_file_dump upc_loop_csv_dumper_62;
    upc_loop_monitor #(34) upc_loop_monitor_62;
    upc_loop_intf#(34) upc_loop_intf_63(clock,reset);
    assign upc_loop_intf_63.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_CS_fsm;
    assign upc_loop_intf_63.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_63.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_63.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_63.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_63.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_63.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_63.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_63.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_63.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_63.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_start;
    assign upc_loop_intf_63.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_ready;
    assign upc_loop_intf_63.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_362_fu_12675.ap_done_int;
    assign upc_loop_intf_63.loop_continue = 1'b1;
    assign upc_loop_intf_63.quit_at_end = 1'b1;
    assign upc_loop_intf_63.finish = finish;
    csv_file_dump upc_loop_csv_dumper_63;
    upc_loop_monitor #(34) upc_loop_monitor_63;
    upc_loop_intf#(34) upc_loop_intf_64(clock,reset);
    assign upc_loop_intf_64.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_CS_fsm;
    assign upc_loop_intf_64.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_64.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_64.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_64.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_64.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_64.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_64.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_64.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_64.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_64.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_start;
    assign upc_loop_intf_64.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_ready;
    assign upc_loop_intf_64.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_363_fu_12717.ap_done_int;
    assign upc_loop_intf_64.loop_continue = 1'b1;
    assign upc_loop_intf_64.quit_at_end = 1'b1;
    assign upc_loop_intf_64.finish = finish;
    csv_file_dump upc_loop_csv_dumper_64;
    upc_loop_monitor #(34) upc_loop_monitor_64;
    upc_loop_intf#(34) upc_loop_intf_65(clock,reset);
    assign upc_loop_intf_65.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_CS_fsm;
    assign upc_loop_intf_65.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_65.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_65.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_65.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_65.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_65.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_65.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_65.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_65.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_65.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_start;
    assign upc_loop_intf_65.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_ready;
    assign upc_loop_intf_65.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_364_fu_12759.ap_done_int;
    assign upc_loop_intf_65.loop_continue = 1'b1;
    assign upc_loop_intf_65.quit_at_end = 1'b1;
    assign upc_loop_intf_65.finish = finish;
    csv_file_dump upc_loop_csv_dumper_65;
    upc_loop_monitor #(34) upc_loop_monitor_65;
    upc_loop_intf#(34) upc_loop_intf_66(clock,reset);
    assign upc_loop_intf_66.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_CS_fsm;
    assign upc_loop_intf_66.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_66.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_66.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_66.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_66.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_66.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_66.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_66.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_66.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_66.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_start;
    assign upc_loop_intf_66.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_ready;
    assign upc_loop_intf_66.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_365_fu_12801.ap_done_int;
    assign upc_loop_intf_66.loop_continue = 1'b1;
    assign upc_loop_intf_66.quit_at_end = 1'b1;
    assign upc_loop_intf_66.finish = finish;
    csv_file_dump upc_loop_csv_dumper_66;
    upc_loop_monitor #(34) upc_loop_monitor_66;
    upc_loop_intf#(34) upc_loop_intf_67(clock,reset);
    assign upc_loop_intf_67.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_CS_fsm;
    assign upc_loop_intf_67.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_67.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_67.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_67.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_67.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_67.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_67.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_67.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_67.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_67.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_start;
    assign upc_loop_intf_67.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_ready;
    assign upc_loop_intf_67.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_366_fu_12843.ap_done_int;
    assign upc_loop_intf_67.loop_continue = 1'b1;
    assign upc_loop_intf_67.quit_at_end = 1'b1;
    assign upc_loop_intf_67.finish = finish;
    csv_file_dump upc_loop_csv_dumper_67;
    upc_loop_monitor #(34) upc_loop_monitor_67;
    upc_loop_intf#(34) upc_loop_intf_68(clock,reset);
    assign upc_loop_intf_68.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_CS_fsm;
    assign upc_loop_intf_68.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_68.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_68.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_68.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_68.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_68.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_68.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_68.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_68.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_68.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_start;
    assign upc_loop_intf_68.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_ready;
    assign upc_loop_intf_68.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_367_fu_12885.ap_done_int;
    assign upc_loop_intf_68.loop_continue = 1'b1;
    assign upc_loop_intf_68.quit_at_end = 1'b1;
    assign upc_loop_intf_68.finish = finish;
    csv_file_dump upc_loop_csv_dumper_68;
    upc_loop_monitor #(34) upc_loop_monitor_68;
    upc_loop_intf#(34) upc_loop_intf_69(clock,reset);
    assign upc_loop_intf_69.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_CS_fsm;
    assign upc_loop_intf_69.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_69.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_69.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_69.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_69.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_69.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_69.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_69.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_69.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_69.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_start;
    assign upc_loop_intf_69.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_ready;
    assign upc_loop_intf_69.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_368_fu_12927.ap_done_int;
    assign upc_loop_intf_69.loop_continue = 1'b1;
    assign upc_loop_intf_69.quit_at_end = 1'b1;
    assign upc_loop_intf_69.finish = finish;
    csv_file_dump upc_loop_csv_dumper_69;
    upc_loop_monitor #(34) upc_loop_monitor_69;
    upc_loop_intf#(34) upc_loop_intf_70(clock,reset);
    assign upc_loop_intf_70.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_CS_fsm;
    assign upc_loop_intf_70.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_70.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_70.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_70.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_70.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_70.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_70.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_70.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_70.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_70.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_start;
    assign upc_loop_intf_70.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_ready;
    assign upc_loop_intf_70.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_369_fu_12969.ap_done_int;
    assign upc_loop_intf_70.loop_continue = 1'b1;
    assign upc_loop_intf_70.quit_at_end = 1'b1;
    assign upc_loop_intf_70.finish = finish;
    csv_file_dump upc_loop_csv_dumper_70;
    upc_loop_monitor #(34) upc_loop_monitor_70;
    upc_loop_intf#(34) upc_loop_intf_71(clock,reset);
    assign upc_loop_intf_71.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_CS_fsm;
    assign upc_loop_intf_71.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_71.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_71.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_71.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_71.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_71.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_71.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_71.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_71.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_71.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_start;
    assign upc_loop_intf_71.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_ready;
    assign upc_loop_intf_71.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_370_fu_13011.ap_done_int;
    assign upc_loop_intf_71.loop_continue = 1'b1;
    assign upc_loop_intf_71.quit_at_end = 1'b1;
    assign upc_loop_intf_71.finish = finish;
    csv_file_dump upc_loop_csv_dumper_71;
    upc_loop_monitor #(34) upc_loop_monitor_71;
    upc_loop_intf#(34) upc_loop_intf_72(clock,reset);
    assign upc_loop_intf_72.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_CS_fsm;
    assign upc_loop_intf_72.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_72.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_72.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_72.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_72.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_72.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_72.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_72.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_72.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_72.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_start;
    assign upc_loop_intf_72.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_ready;
    assign upc_loop_intf_72.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_371_fu_13053.ap_done_int;
    assign upc_loop_intf_72.loop_continue = 1'b1;
    assign upc_loop_intf_72.quit_at_end = 1'b1;
    assign upc_loop_intf_72.finish = finish;
    csv_file_dump upc_loop_csv_dumper_72;
    upc_loop_monitor #(34) upc_loop_monitor_72;
    upc_loop_intf#(34) upc_loop_intf_73(clock,reset);
    assign upc_loop_intf_73.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_CS_fsm;
    assign upc_loop_intf_73.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_73.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_73.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_73.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_73.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_73.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_73.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_73.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_73.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_73.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_start;
    assign upc_loop_intf_73.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_ready;
    assign upc_loop_intf_73.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_372_fu_13095.ap_done_int;
    assign upc_loop_intf_73.loop_continue = 1'b1;
    assign upc_loop_intf_73.quit_at_end = 1'b1;
    assign upc_loop_intf_73.finish = finish;
    csv_file_dump upc_loop_csv_dumper_73;
    upc_loop_monitor #(34) upc_loop_monitor_73;
    upc_loop_intf#(34) upc_loop_intf_74(clock,reset);
    assign upc_loop_intf_74.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_CS_fsm;
    assign upc_loop_intf_74.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_74.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_74.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_74.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_74.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_74.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_74.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_74.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_74.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_74.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_start;
    assign upc_loop_intf_74.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_ready;
    assign upc_loop_intf_74.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_373_fu_13137.ap_done_int;
    assign upc_loop_intf_74.loop_continue = 1'b1;
    assign upc_loop_intf_74.quit_at_end = 1'b1;
    assign upc_loop_intf_74.finish = finish;
    csv_file_dump upc_loop_csv_dumper_74;
    upc_loop_monitor #(34) upc_loop_monitor_74;
    upc_loop_intf#(34) upc_loop_intf_75(clock,reset);
    assign upc_loop_intf_75.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_CS_fsm;
    assign upc_loop_intf_75.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_75.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_75.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_75.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_75.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_75.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_75.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_75.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_75.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_75.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_start;
    assign upc_loop_intf_75.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_ready;
    assign upc_loop_intf_75.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_374_fu_13179.ap_done_int;
    assign upc_loop_intf_75.loop_continue = 1'b1;
    assign upc_loop_intf_75.quit_at_end = 1'b1;
    assign upc_loop_intf_75.finish = finish;
    csv_file_dump upc_loop_csv_dumper_75;
    upc_loop_monitor #(34) upc_loop_monitor_75;
    upc_loop_intf#(34) upc_loop_intf_76(clock,reset);
    assign upc_loop_intf_76.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_CS_fsm;
    assign upc_loop_intf_76.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_76.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_76.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_76.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_76.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_76.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_76.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_76.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_76.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_76.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_start;
    assign upc_loop_intf_76.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_ready;
    assign upc_loop_intf_76.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_375_fu_13221.ap_done_int;
    assign upc_loop_intf_76.loop_continue = 1'b1;
    assign upc_loop_intf_76.quit_at_end = 1'b1;
    assign upc_loop_intf_76.finish = finish;
    csv_file_dump upc_loop_csv_dumper_76;
    upc_loop_monitor #(34) upc_loop_monitor_76;
    upc_loop_intf#(34) upc_loop_intf_77(clock,reset);
    assign upc_loop_intf_77.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_CS_fsm;
    assign upc_loop_intf_77.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_77.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_77.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_77.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_77.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_77.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_77.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_77.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_77.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_77.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_start;
    assign upc_loop_intf_77.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_ready;
    assign upc_loop_intf_77.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_376_fu_13263.ap_done_int;
    assign upc_loop_intf_77.loop_continue = 1'b1;
    assign upc_loop_intf_77.quit_at_end = 1'b1;
    assign upc_loop_intf_77.finish = finish;
    csv_file_dump upc_loop_csv_dumper_77;
    upc_loop_monitor #(34) upc_loop_monitor_77;
    upc_loop_intf#(34) upc_loop_intf_78(clock,reset);
    assign upc_loop_intf_78.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_CS_fsm;
    assign upc_loop_intf_78.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_78.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_78.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_78.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_78.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_78.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_78.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_78.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_78.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_78.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_start;
    assign upc_loop_intf_78.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_ready;
    assign upc_loop_intf_78.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_377_fu_13305.ap_done_int;
    assign upc_loop_intf_78.loop_continue = 1'b1;
    assign upc_loop_intf_78.quit_at_end = 1'b1;
    assign upc_loop_intf_78.finish = finish;
    csv_file_dump upc_loop_csv_dumper_78;
    upc_loop_monitor #(34) upc_loop_monitor_78;
    upc_loop_intf#(34) upc_loop_intf_79(clock,reset);
    assign upc_loop_intf_79.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_CS_fsm;
    assign upc_loop_intf_79.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_79.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_79.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_79.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_79.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_79.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_79.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_79.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_79.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_79.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_start;
    assign upc_loop_intf_79.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_ready;
    assign upc_loop_intf_79.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_378_fu_13347.ap_done_int;
    assign upc_loop_intf_79.loop_continue = 1'b1;
    assign upc_loop_intf_79.quit_at_end = 1'b1;
    assign upc_loop_intf_79.finish = finish;
    csv_file_dump upc_loop_csv_dumper_79;
    upc_loop_monitor #(34) upc_loop_monitor_79;
    upc_loop_intf#(34) upc_loop_intf_80(clock,reset);
    assign upc_loop_intf_80.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_CS_fsm;
    assign upc_loop_intf_80.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_80.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_80.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_80.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_80.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_80.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_80.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_80.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_80.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_80.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_start;
    assign upc_loop_intf_80.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_ready;
    assign upc_loop_intf_80.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_379_fu_13389.ap_done_int;
    assign upc_loop_intf_80.loop_continue = 1'b1;
    assign upc_loop_intf_80.quit_at_end = 1'b1;
    assign upc_loop_intf_80.finish = finish;
    csv_file_dump upc_loop_csv_dumper_80;
    upc_loop_monitor #(34) upc_loop_monitor_80;
    upc_loop_intf#(34) upc_loop_intf_81(clock,reset);
    assign upc_loop_intf_81.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_CS_fsm;
    assign upc_loop_intf_81.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_81.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_81.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_81.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_81.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_81.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_81.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_81.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_81.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_81.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_start;
    assign upc_loop_intf_81.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_ready;
    assign upc_loop_intf_81.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_380_fu_13431.ap_done_int;
    assign upc_loop_intf_81.loop_continue = 1'b1;
    assign upc_loop_intf_81.quit_at_end = 1'b1;
    assign upc_loop_intf_81.finish = finish;
    csv_file_dump upc_loop_csv_dumper_81;
    upc_loop_monitor #(34) upc_loop_monitor_81;
    upc_loop_intf#(34) upc_loop_intf_82(clock,reset);
    assign upc_loop_intf_82.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_CS_fsm;
    assign upc_loop_intf_82.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_82.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_82.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_82.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_82.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_82.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_82.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_82.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_82.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_82.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_start;
    assign upc_loop_intf_82.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_ready;
    assign upc_loop_intf_82.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_381_fu_13473.ap_done_int;
    assign upc_loop_intf_82.loop_continue = 1'b1;
    assign upc_loop_intf_82.quit_at_end = 1'b1;
    assign upc_loop_intf_82.finish = finish;
    csv_file_dump upc_loop_csv_dumper_82;
    upc_loop_monitor #(34) upc_loop_monitor_82;
    upc_loop_intf#(34) upc_loop_intf_83(clock,reset);
    assign upc_loop_intf_83.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_CS_fsm;
    assign upc_loop_intf_83.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_83.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_83.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_83.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_83.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_83.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_83.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_83.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_83.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_83.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_start;
    assign upc_loop_intf_83.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_ready;
    assign upc_loop_intf_83.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_382_fu_13515.ap_done_int;
    assign upc_loop_intf_83.loop_continue = 1'b1;
    assign upc_loop_intf_83.quit_at_end = 1'b1;
    assign upc_loop_intf_83.finish = finish;
    csv_file_dump upc_loop_csv_dumper_83;
    upc_loop_monitor #(34) upc_loop_monitor_83;
    upc_loop_intf#(34) upc_loop_intf_84(clock,reset);
    assign upc_loop_intf_84.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_CS_fsm;
    assign upc_loop_intf_84.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_84.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_84.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_84.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_84.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_84.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_84.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_84.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_84.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_84.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_start;
    assign upc_loop_intf_84.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_ready;
    assign upc_loop_intf_84.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_383_fu_13557.ap_done_int;
    assign upc_loop_intf_84.loop_continue = 1'b1;
    assign upc_loop_intf_84.quit_at_end = 1'b1;
    assign upc_loop_intf_84.finish = finish;
    csv_file_dump upc_loop_csv_dumper_84;
    upc_loop_monitor #(34) upc_loop_monitor_84;
    upc_loop_intf#(34) upc_loop_intf_85(clock,reset);
    assign upc_loop_intf_85.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_CS_fsm;
    assign upc_loop_intf_85.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_85.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_85.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_85.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_85.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_85.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_85.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_85.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_85.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_85.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_start;
    assign upc_loop_intf_85.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_ready;
    assign upc_loop_intf_85.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_384_fu_13599.ap_done_int;
    assign upc_loop_intf_85.loop_continue = 1'b1;
    assign upc_loop_intf_85.quit_at_end = 1'b1;
    assign upc_loop_intf_85.finish = finish;
    csv_file_dump upc_loop_csv_dumper_85;
    upc_loop_monitor #(34) upc_loop_monitor_85;
    upc_loop_intf#(34) upc_loop_intf_86(clock,reset);
    assign upc_loop_intf_86.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_CS_fsm;
    assign upc_loop_intf_86.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_86.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_86.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_86.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_86.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_86.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_86.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_86.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_86.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_86.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_start;
    assign upc_loop_intf_86.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_ready;
    assign upc_loop_intf_86.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_385_fu_13641.ap_done_int;
    assign upc_loop_intf_86.loop_continue = 1'b1;
    assign upc_loop_intf_86.quit_at_end = 1'b1;
    assign upc_loop_intf_86.finish = finish;
    csv_file_dump upc_loop_csv_dumper_86;
    upc_loop_monitor #(34) upc_loop_monitor_86;
    upc_loop_intf#(34) upc_loop_intf_87(clock,reset);
    assign upc_loop_intf_87.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_CS_fsm;
    assign upc_loop_intf_87.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_87.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_87.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_87.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_87.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_87.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_87.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_87.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_87.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_87.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_start;
    assign upc_loop_intf_87.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_ready;
    assign upc_loop_intf_87.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_386_fu_13683.ap_done_int;
    assign upc_loop_intf_87.loop_continue = 1'b1;
    assign upc_loop_intf_87.quit_at_end = 1'b1;
    assign upc_loop_intf_87.finish = finish;
    csv_file_dump upc_loop_csv_dumper_87;
    upc_loop_monitor #(34) upc_loop_monitor_87;
    upc_loop_intf#(34) upc_loop_intf_88(clock,reset);
    assign upc_loop_intf_88.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_CS_fsm;
    assign upc_loop_intf_88.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_88.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_88.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_88.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_88.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_88.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_88.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_88.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_88.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_88.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_start;
    assign upc_loop_intf_88.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_ready;
    assign upc_loop_intf_88.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_387_fu_13725.ap_done_int;
    assign upc_loop_intf_88.loop_continue = 1'b1;
    assign upc_loop_intf_88.quit_at_end = 1'b1;
    assign upc_loop_intf_88.finish = finish;
    csv_file_dump upc_loop_csv_dumper_88;
    upc_loop_monitor #(34) upc_loop_monitor_88;
    upc_loop_intf#(34) upc_loop_intf_89(clock,reset);
    assign upc_loop_intf_89.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_CS_fsm;
    assign upc_loop_intf_89.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_89.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_89.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_89.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_89.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_89.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_89.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_89.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_89.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_89.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_start;
    assign upc_loop_intf_89.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_ready;
    assign upc_loop_intf_89.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_388_fu_13767.ap_done_int;
    assign upc_loop_intf_89.loop_continue = 1'b1;
    assign upc_loop_intf_89.quit_at_end = 1'b1;
    assign upc_loop_intf_89.finish = finish;
    csv_file_dump upc_loop_csv_dumper_89;
    upc_loop_monitor #(34) upc_loop_monitor_89;
    upc_loop_intf#(34) upc_loop_intf_90(clock,reset);
    assign upc_loop_intf_90.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_CS_fsm;
    assign upc_loop_intf_90.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_90.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_90.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_90.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_90.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_90.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_90.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_90.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_90.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_90.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_start;
    assign upc_loop_intf_90.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_ready;
    assign upc_loop_intf_90.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_389_fu_13809.ap_done_int;
    assign upc_loop_intf_90.loop_continue = 1'b1;
    assign upc_loop_intf_90.quit_at_end = 1'b1;
    assign upc_loop_intf_90.finish = finish;
    csv_file_dump upc_loop_csv_dumper_90;
    upc_loop_monitor #(34) upc_loop_monitor_90;
    upc_loop_intf#(34) upc_loop_intf_91(clock,reset);
    assign upc_loop_intf_91.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_CS_fsm;
    assign upc_loop_intf_91.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_91.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_91.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_91.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_91.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_91.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_91.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_91.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_91.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_91.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_start;
    assign upc_loop_intf_91.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_ready;
    assign upc_loop_intf_91.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_390_fu_13851.ap_done_int;
    assign upc_loop_intf_91.loop_continue = 1'b1;
    assign upc_loop_intf_91.quit_at_end = 1'b1;
    assign upc_loop_intf_91.finish = finish;
    csv_file_dump upc_loop_csv_dumper_91;
    upc_loop_monitor #(34) upc_loop_monitor_91;
    upc_loop_intf#(34) upc_loop_intf_92(clock,reset);
    assign upc_loop_intf_92.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_CS_fsm;
    assign upc_loop_intf_92.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_92.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_92.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_92.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_92.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_92.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_92.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_92.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_92.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_92.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_start;
    assign upc_loop_intf_92.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_ready;
    assign upc_loop_intf_92.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_391_fu_13893.ap_done_int;
    assign upc_loop_intf_92.loop_continue = 1'b1;
    assign upc_loop_intf_92.quit_at_end = 1'b1;
    assign upc_loop_intf_92.finish = finish;
    csv_file_dump upc_loop_csv_dumper_92;
    upc_loop_monitor #(34) upc_loop_monitor_92;
    upc_loop_intf#(34) upc_loop_intf_93(clock,reset);
    assign upc_loop_intf_93.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_CS_fsm;
    assign upc_loop_intf_93.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_93.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_93.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_93.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_93.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_93.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_93.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_93.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_93.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_93.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_start;
    assign upc_loop_intf_93.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_ready;
    assign upc_loop_intf_93.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_392_fu_13935.ap_done_int;
    assign upc_loop_intf_93.loop_continue = 1'b1;
    assign upc_loop_intf_93.quit_at_end = 1'b1;
    assign upc_loop_intf_93.finish = finish;
    csv_file_dump upc_loop_csv_dumper_93;
    upc_loop_monitor #(34) upc_loop_monitor_93;
    upc_loop_intf#(34) upc_loop_intf_94(clock,reset);
    assign upc_loop_intf_94.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_CS_fsm;
    assign upc_loop_intf_94.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_94.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_94.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_94.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_94.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_94.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_94.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_94.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_94.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_94.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_start;
    assign upc_loop_intf_94.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_ready;
    assign upc_loop_intf_94.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_393_fu_13977.ap_done_int;
    assign upc_loop_intf_94.loop_continue = 1'b1;
    assign upc_loop_intf_94.quit_at_end = 1'b1;
    assign upc_loop_intf_94.finish = finish;
    csv_file_dump upc_loop_csv_dumper_94;
    upc_loop_monitor #(34) upc_loop_monitor_94;
    upc_loop_intf#(34) upc_loop_intf_95(clock,reset);
    assign upc_loop_intf_95.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_CS_fsm;
    assign upc_loop_intf_95.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_95.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_95.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_95.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_95.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_95.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_95.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_95.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_95.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_95.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_start;
    assign upc_loop_intf_95.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_ready;
    assign upc_loop_intf_95.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_394_fu_14019.ap_done_int;
    assign upc_loop_intf_95.loop_continue = 1'b1;
    assign upc_loop_intf_95.quit_at_end = 1'b1;
    assign upc_loop_intf_95.finish = finish;
    csv_file_dump upc_loop_csv_dumper_95;
    upc_loop_monitor #(34) upc_loop_monitor_95;
    upc_loop_intf#(34) upc_loop_intf_96(clock,reset);
    assign upc_loop_intf_96.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_CS_fsm;
    assign upc_loop_intf_96.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_96.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_96.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_96.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_96.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_96.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_96.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_96.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_96.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_96.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_start;
    assign upc_loop_intf_96.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_ready;
    assign upc_loop_intf_96.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_395_fu_14061.ap_done_int;
    assign upc_loop_intf_96.loop_continue = 1'b1;
    assign upc_loop_intf_96.quit_at_end = 1'b1;
    assign upc_loop_intf_96.finish = finish;
    csv_file_dump upc_loop_csv_dumper_96;
    upc_loop_monitor #(34) upc_loop_monitor_96;
    upc_loop_intf#(34) upc_loop_intf_97(clock,reset);
    assign upc_loop_intf_97.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_CS_fsm;
    assign upc_loop_intf_97.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_97.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_97.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_97.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_97.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_97.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_97.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_97.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_97.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_97.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_start;
    assign upc_loop_intf_97.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_ready;
    assign upc_loop_intf_97.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_396_fu_14103.ap_done_int;
    assign upc_loop_intf_97.loop_continue = 1'b1;
    assign upc_loop_intf_97.quit_at_end = 1'b1;
    assign upc_loop_intf_97.finish = finish;
    csv_file_dump upc_loop_csv_dumper_97;
    upc_loop_monitor #(34) upc_loop_monitor_97;
    upc_loop_intf#(34) upc_loop_intf_98(clock,reset);
    assign upc_loop_intf_98.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_CS_fsm;
    assign upc_loop_intf_98.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_98.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_98.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_98.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_98.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_98.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_98.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_98.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_98.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_98.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_start;
    assign upc_loop_intf_98.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_ready;
    assign upc_loop_intf_98.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_397_fu_14145.ap_done_int;
    assign upc_loop_intf_98.loop_continue = 1'b1;
    assign upc_loop_intf_98.quit_at_end = 1'b1;
    assign upc_loop_intf_98.finish = finish;
    csv_file_dump upc_loop_csv_dumper_98;
    upc_loop_monitor #(34) upc_loop_monitor_98;
    upc_loop_intf#(34) upc_loop_intf_99(clock,reset);
    assign upc_loop_intf_99.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_CS_fsm;
    assign upc_loop_intf_99.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_99.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_99.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_99.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_99.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_99.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_99.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_99.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_99.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_99.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_start;
    assign upc_loop_intf_99.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_ready;
    assign upc_loop_intf_99.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_398_fu_14187.ap_done_int;
    assign upc_loop_intf_99.loop_continue = 1'b1;
    assign upc_loop_intf_99.quit_at_end = 1'b1;
    assign upc_loop_intf_99.finish = finish;
    csv_file_dump upc_loop_csv_dumper_99;
    upc_loop_monitor #(34) upc_loop_monitor_99;
    upc_loop_intf#(34) upc_loop_intf_100(clock,reset);
    assign upc_loop_intf_100.cur_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_CS_fsm;
    assign upc_loop_intf_100.iter_start_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_100.iter_end_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_100.quit_state = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_ST_fsm_pp0_stage10;
    assign upc_loop_intf_100.iter_start_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_100.iter_end_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_100.quit_block = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_block_pp0_stage10_subdone;
    assign upc_loop_intf_100.iter_start_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_100.iter_end_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_100.quit_enable = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_100.loop_start = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_start;
    assign upc_loop_intf_100.loop_ready = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_ready;
    assign upc_loop_intf_100.loop_done = AESL_inst_SABR.grp_SABR_Pipeline_VITIS_LOOP_31_399_fu_14229.ap_done_int;
    assign upc_loop_intf_100.loop_continue = 1'b1;
    assign upc_loop_intf_100.quit_at_end = 1'b1;
    assign upc_loop_intf_100.finish = finish;
    csv_file_dump upc_loop_csv_dumper_100;
    upc_loop_monitor #(34) upc_loop_monitor_100;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);
    mstatus_csv_dumper_68 = new("./module_status68.csv");
    module_monitor_68 = new(module_intf_68,mstatus_csv_dumper_68);
    mstatus_csv_dumper_69 = new("./module_status69.csv");
    module_monitor_69 = new(module_intf_69,mstatus_csv_dumper_69);
    mstatus_csv_dumper_70 = new("./module_status70.csv");
    module_monitor_70 = new(module_intf_70,mstatus_csv_dumper_70);
    mstatus_csv_dumper_71 = new("./module_status71.csv");
    module_monitor_71 = new(module_intf_71,mstatus_csv_dumper_71);
    mstatus_csv_dumper_72 = new("./module_status72.csv");
    module_monitor_72 = new(module_intf_72,mstatus_csv_dumper_72);
    mstatus_csv_dumper_73 = new("./module_status73.csv");
    module_monitor_73 = new(module_intf_73,mstatus_csv_dumper_73);
    mstatus_csv_dumper_74 = new("./module_status74.csv");
    module_monitor_74 = new(module_intf_74,mstatus_csv_dumper_74);
    mstatus_csv_dumper_75 = new("./module_status75.csv");
    module_monitor_75 = new(module_intf_75,mstatus_csv_dumper_75);
    mstatus_csv_dumper_76 = new("./module_status76.csv");
    module_monitor_76 = new(module_intf_76,mstatus_csv_dumper_76);
    mstatus_csv_dumper_77 = new("./module_status77.csv");
    module_monitor_77 = new(module_intf_77,mstatus_csv_dumper_77);
    mstatus_csv_dumper_78 = new("./module_status78.csv");
    module_monitor_78 = new(module_intf_78,mstatus_csv_dumper_78);
    mstatus_csv_dumper_79 = new("./module_status79.csv");
    module_monitor_79 = new(module_intf_79,mstatus_csv_dumper_79);
    mstatus_csv_dumper_80 = new("./module_status80.csv");
    module_monitor_80 = new(module_intf_80,mstatus_csv_dumper_80);
    mstatus_csv_dumper_81 = new("./module_status81.csv");
    module_monitor_81 = new(module_intf_81,mstatus_csv_dumper_81);
    mstatus_csv_dumper_82 = new("./module_status82.csv");
    module_monitor_82 = new(module_intf_82,mstatus_csv_dumper_82);
    mstatus_csv_dumper_83 = new("./module_status83.csv");
    module_monitor_83 = new(module_intf_83,mstatus_csv_dumper_83);
    mstatus_csv_dumper_84 = new("./module_status84.csv");
    module_monitor_84 = new(module_intf_84,mstatus_csv_dumper_84);
    mstatus_csv_dumper_85 = new("./module_status85.csv");
    module_monitor_85 = new(module_intf_85,mstatus_csv_dumper_85);
    mstatus_csv_dumper_86 = new("./module_status86.csv");
    module_monitor_86 = new(module_intf_86,mstatus_csv_dumper_86);
    mstatus_csv_dumper_87 = new("./module_status87.csv");
    module_monitor_87 = new(module_intf_87,mstatus_csv_dumper_87);
    mstatus_csv_dumper_88 = new("./module_status88.csv");
    module_monitor_88 = new(module_intf_88,mstatus_csv_dumper_88);
    mstatus_csv_dumper_89 = new("./module_status89.csv");
    module_monitor_89 = new(module_intf_89,mstatus_csv_dumper_89);
    mstatus_csv_dumper_90 = new("./module_status90.csv");
    module_monitor_90 = new(module_intf_90,mstatus_csv_dumper_90);
    mstatus_csv_dumper_91 = new("./module_status91.csv");
    module_monitor_91 = new(module_intf_91,mstatus_csv_dumper_91);
    mstatus_csv_dumper_92 = new("./module_status92.csv");
    module_monitor_92 = new(module_intf_92,mstatus_csv_dumper_92);
    mstatus_csv_dumper_93 = new("./module_status93.csv");
    module_monitor_93 = new(module_intf_93,mstatus_csv_dumper_93);
    mstatus_csv_dumper_94 = new("./module_status94.csv");
    module_monitor_94 = new(module_intf_94,mstatus_csv_dumper_94);
    mstatus_csv_dumper_95 = new("./module_status95.csv");
    module_monitor_95 = new(module_intf_95,mstatus_csv_dumper_95);
    mstatus_csv_dumper_96 = new("./module_status96.csv");
    module_monitor_96 = new(module_intf_96,mstatus_csv_dumper_96);
    mstatus_csv_dumper_97 = new("./module_status97.csv");
    module_monitor_97 = new(module_intf_97,mstatus_csv_dumper_97);
    mstatus_csv_dumper_98 = new("./module_status98.csv");
    module_monitor_98 = new(module_intf_98,mstatus_csv_dumper_98);
    mstatus_csv_dumper_99 = new("./module_status99.csv");
    module_monitor_99 = new(module_intf_99,mstatus_csv_dumper_99);
    mstatus_csv_dumper_100 = new("./module_status100.csv");
    module_monitor_100 = new(module_intf_100,mstatus_csv_dumper_100);
    mstatus_csv_dumper_101 = new("./module_status101.csv");
    module_monitor_101 = new(module_intf_101,mstatus_csv_dumper_101);
    mstatus_csv_dumper_102 = new("./module_status102.csv");
    module_monitor_102 = new(module_intf_102,mstatus_csv_dumper_102);




    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);
    upc_loop_csv_dumper_24 = new("./upc_loop_status24.csv");
    upc_loop_monitor_24 = new(upc_loop_intf_24,upc_loop_csv_dumper_24);
    upc_loop_csv_dumper_25 = new("./upc_loop_status25.csv");
    upc_loop_monitor_25 = new(upc_loop_intf_25,upc_loop_csv_dumper_25);
    upc_loop_csv_dumper_26 = new("./upc_loop_status26.csv");
    upc_loop_monitor_26 = new(upc_loop_intf_26,upc_loop_csv_dumper_26);
    upc_loop_csv_dumper_27 = new("./upc_loop_status27.csv");
    upc_loop_monitor_27 = new(upc_loop_intf_27,upc_loop_csv_dumper_27);
    upc_loop_csv_dumper_28 = new("./upc_loop_status28.csv");
    upc_loop_monitor_28 = new(upc_loop_intf_28,upc_loop_csv_dumper_28);
    upc_loop_csv_dumper_29 = new("./upc_loop_status29.csv");
    upc_loop_monitor_29 = new(upc_loop_intf_29,upc_loop_csv_dumper_29);
    upc_loop_csv_dumper_30 = new("./upc_loop_status30.csv");
    upc_loop_monitor_30 = new(upc_loop_intf_30,upc_loop_csv_dumper_30);
    upc_loop_csv_dumper_31 = new("./upc_loop_status31.csv");
    upc_loop_monitor_31 = new(upc_loop_intf_31,upc_loop_csv_dumper_31);
    upc_loop_csv_dumper_32 = new("./upc_loop_status32.csv");
    upc_loop_monitor_32 = new(upc_loop_intf_32,upc_loop_csv_dumper_32);
    upc_loop_csv_dumper_33 = new("./upc_loop_status33.csv");
    upc_loop_monitor_33 = new(upc_loop_intf_33,upc_loop_csv_dumper_33);
    upc_loop_csv_dumper_34 = new("./upc_loop_status34.csv");
    upc_loop_monitor_34 = new(upc_loop_intf_34,upc_loop_csv_dumper_34);
    upc_loop_csv_dumper_35 = new("./upc_loop_status35.csv");
    upc_loop_monitor_35 = new(upc_loop_intf_35,upc_loop_csv_dumper_35);
    upc_loop_csv_dumper_36 = new("./upc_loop_status36.csv");
    upc_loop_monitor_36 = new(upc_loop_intf_36,upc_loop_csv_dumper_36);
    upc_loop_csv_dumper_37 = new("./upc_loop_status37.csv");
    upc_loop_monitor_37 = new(upc_loop_intf_37,upc_loop_csv_dumper_37);
    upc_loop_csv_dumper_38 = new("./upc_loop_status38.csv");
    upc_loop_monitor_38 = new(upc_loop_intf_38,upc_loop_csv_dumper_38);
    upc_loop_csv_dumper_39 = new("./upc_loop_status39.csv");
    upc_loop_monitor_39 = new(upc_loop_intf_39,upc_loop_csv_dumper_39);
    upc_loop_csv_dumper_40 = new("./upc_loop_status40.csv");
    upc_loop_monitor_40 = new(upc_loop_intf_40,upc_loop_csv_dumper_40);
    upc_loop_csv_dumper_41 = new("./upc_loop_status41.csv");
    upc_loop_monitor_41 = new(upc_loop_intf_41,upc_loop_csv_dumper_41);
    upc_loop_csv_dumper_42 = new("./upc_loop_status42.csv");
    upc_loop_monitor_42 = new(upc_loop_intf_42,upc_loop_csv_dumper_42);
    upc_loop_csv_dumper_43 = new("./upc_loop_status43.csv");
    upc_loop_monitor_43 = new(upc_loop_intf_43,upc_loop_csv_dumper_43);
    upc_loop_csv_dumper_44 = new("./upc_loop_status44.csv");
    upc_loop_monitor_44 = new(upc_loop_intf_44,upc_loop_csv_dumper_44);
    upc_loop_csv_dumper_45 = new("./upc_loop_status45.csv");
    upc_loop_monitor_45 = new(upc_loop_intf_45,upc_loop_csv_dumper_45);
    upc_loop_csv_dumper_46 = new("./upc_loop_status46.csv");
    upc_loop_monitor_46 = new(upc_loop_intf_46,upc_loop_csv_dumper_46);
    upc_loop_csv_dumper_47 = new("./upc_loop_status47.csv");
    upc_loop_monitor_47 = new(upc_loop_intf_47,upc_loop_csv_dumper_47);
    upc_loop_csv_dumper_48 = new("./upc_loop_status48.csv");
    upc_loop_monitor_48 = new(upc_loop_intf_48,upc_loop_csv_dumper_48);
    upc_loop_csv_dumper_49 = new("./upc_loop_status49.csv");
    upc_loop_monitor_49 = new(upc_loop_intf_49,upc_loop_csv_dumper_49);
    upc_loop_csv_dumper_50 = new("./upc_loop_status50.csv");
    upc_loop_monitor_50 = new(upc_loop_intf_50,upc_loop_csv_dumper_50);
    upc_loop_csv_dumper_51 = new("./upc_loop_status51.csv");
    upc_loop_monitor_51 = new(upc_loop_intf_51,upc_loop_csv_dumper_51);
    upc_loop_csv_dumper_52 = new("./upc_loop_status52.csv");
    upc_loop_monitor_52 = new(upc_loop_intf_52,upc_loop_csv_dumper_52);
    upc_loop_csv_dumper_53 = new("./upc_loop_status53.csv");
    upc_loop_monitor_53 = new(upc_loop_intf_53,upc_loop_csv_dumper_53);
    upc_loop_csv_dumper_54 = new("./upc_loop_status54.csv");
    upc_loop_monitor_54 = new(upc_loop_intf_54,upc_loop_csv_dumper_54);
    upc_loop_csv_dumper_55 = new("./upc_loop_status55.csv");
    upc_loop_monitor_55 = new(upc_loop_intf_55,upc_loop_csv_dumper_55);
    upc_loop_csv_dumper_56 = new("./upc_loop_status56.csv");
    upc_loop_monitor_56 = new(upc_loop_intf_56,upc_loop_csv_dumper_56);
    upc_loop_csv_dumper_57 = new("./upc_loop_status57.csv");
    upc_loop_monitor_57 = new(upc_loop_intf_57,upc_loop_csv_dumper_57);
    upc_loop_csv_dumper_58 = new("./upc_loop_status58.csv");
    upc_loop_monitor_58 = new(upc_loop_intf_58,upc_loop_csv_dumper_58);
    upc_loop_csv_dumper_59 = new("./upc_loop_status59.csv");
    upc_loop_monitor_59 = new(upc_loop_intf_59,upc_loop_csv_dumper_59);
    upc_loop_csv_dumper_60 = new("./upc_loop_status60.csv");
    upc_loop_monitor_60 = new(upc_loop_intf_60,upc_loop_csv_dumper_60);
    upc_loop_csv_dumper_61 = new("./upc_loop_status61.csv");
    upc_loop_monitor_61 = new(upc_loop_intf_61,upc_loop_csv_dumper_61);
    upc_loop_csv_dumper_62 = new("./upc_loop_status62.csv");
    upc_loop_monitor_62 = new(upc_loop_intf_62,upc_loop_csv_dumper_62);
    upc_loop_csv_dumper_63 = new("./upc_loop_status63.csv");
    upc_loop_monitor_63 = new(upc_loop_intf_63,upc_loop_csv_dumper_63);
    upc_loop_csv_dumper_64 = new("./upc_loop_status64.csv");
    upc_loop_monitor_64 = new(upc_loop_intf_64,upc_loop_csv_dumper_64);
    upc_loop_csv_dumper_65 = new("./upc_loop_status65.csv");
    upc_loop_monitor_65 = new(upc_loop_intf_65,upc_loop_csv_dumper_65);
    upc_loop_csv_dumper_66 = new("./upc_loop_status66.csv");
    upc_loop_monitor_66 = new(upc_loop_intf_66,upc_loop_csv_dumper_66);
    upc_loop_csv_dumper_67 = new("./upc_loop_status67.csv");
    upc_loop_monitor_67 = new(upc_loop_intf_67,upc_loop_csv_dumper_67);
    upc_loop_csv_dumper_68 = new("./upc_loop_status68.csv");
    upc_loop_monitor_68 = new(upc_loop_intf_68,upc_loop_csv_dumper_68);
    upc_loop_csv_dumper_69 = new("./upc_loop_status69.csv");
    upc_loop_monitor_69 = new(upc_loop_intf_69,upc_loop_csv_dumper_69);
    upc_loop_csv_dumper_70 = new("./upc_loop_status70.csv");
    upc_loop_monitor_70 = new(upc_loop_intf_70,upc_loop_csv_dumper_70);
    upc_loop_csv_dumper_71 = new("./upc_loop_status71.csv");
    upc_loop_monitor_71 = new(upc_loop_intf_71,upc_loop_csv_dumper_71);
    upc_loop_csv_dumper_72 = new("./upc_loop_status72.csv");
    upc_loop_monitor_72 = new(upc_loop_intf_72,upc_loop_csv_dumper_72);
    upc_loop_csv_dumper_73 = new("./upc_loop_status73.csv");
    upc_loop_monitor_73 = new(upc_loop_intf_73,upc_loop_csv_dumper_73);
    upc_loop_csv_dumper_74 = new("./upc_loop_status74.csv");
    upc_loop_monitor_74 = new(upc_loop_intf_74,upc_loop_csv_dumper_74);
    upc_loop_csv_dumper_75 = new("./upc_loop_status75.csv");
    upc_loop_monitor_75 = new(upc_loop_intf_75,upc_loop_csv_dumper_75);
    upc_loop_csv_dumper_76 = new("./upc_loop_status76.csv");
    upc_loop_monitor_76 = new(upc_loop_intf_76,upc_loop_csv_dumper_76);
    upc_loop_csv_dumper_77 = new("./upc_loop_status77.csv");
    upc_loop_monitor_77 = new(upc_loop_intf_77,upc_loop_csv_dumper_77);
    upc_loop_csv_dumper_78 = new("./upc_loop_status78.csv");
    upc_loop_monitor_78 = new(upc_loop_intf_78,upc_loop_csv_dumper_78);
    upc_loop_csv_dumper_79 = new("./upc_loop_status79.csv");
    upc_loop_monitor_79 = new(upc_loop_intf_79,upc_loop_csv_dumper_79);
    upc_loop_csv_dumper_80 = new("./upc_loop_status80.csv");
    upc_loop_monitor_80 = new(upc_loop_intf_80,upc_loop_csv_dumper_80);
    upc_loop_csv_dumper_81 = new("./upc_loop_status81.csv");
    upc_loop_monitor_81 = new(upc_loop_intf_81,upc_loop_csv_dumper_81);
    upc_loop_csv_dumper_82 = new("./upc_loop_status82.csv");
    upc_loop_monitor_82 = new(upc_loop_intf_82,upc_loop_csv_dumper_82);
    upc_loop_csv_dumper_83 = new("./upc_loop_status83.csv");
    upc_loop_monitor_83 = new(upc_loop_intf_83,upc_loop_csv_dumper_83);
    upc_loop_csv_dumper_84 = new("./upc_loop_status84.csv");
    upc_loop_monitor_84 = new(upc_loop_intf_84,upc_loop_csv_dumper_84);
    upc_loop_csv_dumper_85 = new("./upc_loop_status85.csv");
    upc_loop_monitor_85 = new(upc_loop_intf_85,upc_loop_csv_dumper_85);
    upc_loop_csv_dumper_86 = new("./upc_loop_status86.csv");
    upc_loop_monitor_86 = new(upc_loop_intf_86,upc_loop_csv_dumper_86);
    upc_loop_csv_dumper_87 = new("./upc_loop_status87.csv");
    upc_loop_monitor_87 = new(upc_loop_intf_87,upc_loop_csv_dumper_87);
    upc_loop_csv_dumper_88 = new("./upc_loop_status88.csv");
    upc_loop_monitor_88 = new(upc_loop_intf_88,upc_loop_csv_dumper_88);
    upc_loop_csv_dumper_89 = new("./upc_loop_status89.csv");
    upc_loop_monitor_89 = new(upc_loop_intf_89,upc_loop_csv_dumper_89);
    upc_loop_csv_dumper_90 = new("./upc_loop_status90.csv");
    upc_loop_monitor_90 = new(upc_loop_intf_90,upc_loop_csv_dumper_90);
    upc_loop_csv_dumper_91 = new("./upc_loop_status91.csv");
    upc_loop_monitor_91 = new(upc_loop_intf_91,upc_loop_csv_dumper_91);
    upc_loop_csv_dumper_92 = new("./upc_loop_status92.csv");
    upc_loop_monitor_92 = new(upc_loop_intf_92,upc_loop_csv_dumper_92);
    upc_loop_csv_dumper_93 = new("./upc_loop_status93.csv");
    upc_loop_monitor_93 = new(upc_loop_intf_93,upc_loop_csv_dumper_93);
    upc_loop_csv_dumper_94 = new("./upc_loop_status94.csv");
    upc_loop_monitor_94 = new(upc_loop_intf_94,upc_loop_csv_dumper_94);
    upc_loop_csv_dumper_95 = new("./upc_loop_status95.csv");
    upc_loop_monitor_95 = new(upc_loop_intf_95,upc_loop_csv_dumper_95);
    upc_loop_csv_dumper_96 = new("./upc_loop_status96.csv");
    upc_loop_monitor_96 = new(upc_loop_intf_96,upc_loop_csv_dumper_96);
    upc_loop_csv_dumper_97 = new("./upc_loop_status97.csv");
    upc_loop_monitor_97 = new(upc_loop_intf_97,upc_loop_csv_dumper_97);
    upc_loop_csv_dumper_98 = new("./upc_loop_status98.csv");
    upc_loop_monitor_98 = new(upc_loop_intf_98,upc_loop_csv_dumper_98);
    upc_loop_csv_dumper_99 = new("./upc_loop_status99.csv");
    upc_loop_monitor_99 = new(upc_loop_intf_99,upc_loop_csv_dumper_99);
    upc_loop_csv_dumper_100 = new("./upc_loop_status100.csv");
    upc_loop_monitor_100 = new(upc_loop_intf_100,upc_loop_csv_dumper_100);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(module_monitor_68);
    sample_manager_inst.add_one_monitor(module_monitor_69);
    sample_manager_inst.add_one_monitor(module_monitor_70);
    sample_manager_inst.add_one_monitor(module_monitor_71);
    sample_manager_inst.add_one_monitor(module_monitor_72);
    sample_manager_inst.add_one_monitor(module_monitor_73);
    sample_manager_inst.add_one_monitor(module_monitor_74);
    sample_manager_inst.add_one_monitor(module_monitor_75);
    sample_manager_inst.add_one_monitor(module_monitor_76);
    sample_manager_inst.add_one_monitor(module_monitor_77);
    sample_manager_inst.add_one_monitor(module_monitor_78);
    sample_manager_inst.add_one_monitor(module_monitor_79);
    sample_manager_inst.add_one_monitor(module_monitor_80);
    sample_manager_inst.add_one_monitor(module_monitor_81);
    sample_manager_inst.add_one_monitor(module_monitor_82);
    sample_manager_inst.add_one_monitor(module_monitor_83);
    sample_manager_inst.add_one_monitor(module_monitor_84);
    sample_manager_inst.add_one_monitor(module_monitor_85);
    sample_manager_inst.add_one_monitor(module_monitor_86);
    sample_manager_inst.add_one_monitor(module_monitor_87);
    sample_manager_inst.add_one_monitor(module_monitor_88);
    sample_manager_inst.add_one_monitor(module_monitor_89);
    sample_manager_inst.add_one_monitor(module_monitor_90);
    sample_manager_inst.add_one_monitor(module_monitor_91);
    sample_manager_inst.add_one_monitor(module_monitor_92);
    sample_manager_inst.add_one_monitor(module_monitor_93);
    sample_manager_inst.add_one_monitor(module_monitor_94);
    sample_manager_inst.add_one_monitor(module_monitor_95);
    sample_manager_inst.add_one_monitor(module_monitor_96);
    sample_manager_inst.add_one_monitor(module_monitor_97);
    sample_manager_inst.add_one_monitor(module_monitor_98);
    sample_manager_inst.add_one_monitor(module_monitor_99);
    sample_manager_inst.add_one_monitor(module_monitor_100);
    sample_manager_inst.add_one_monitor(module_monitor_101);
    sample_manager_inst.add_one_monitor(module_monitor_102);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_24);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_26);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_27);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_28);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_29);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_30);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_31);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_32);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_33);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_34);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_35);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_36);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_37);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_38);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_39);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_40);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_41);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_42);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_43);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_44);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_45);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_46);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_47);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_48);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_49);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_50);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_51);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_52);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_53);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_54);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_55);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_56);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_57);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_58);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_59);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_60);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_61);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_62);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_63);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_64);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_65);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_66);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_67);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_68);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_69);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_70);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_71);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_72);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_73);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_74);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_75);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_76);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_77);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_78);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_79);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_80);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_81);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_82);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_83);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_84);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_85);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_86);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_87);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_88);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_89);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_90);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_91);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_92);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_93);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_94);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_95);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_96);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_97);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_98);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_99);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_100);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
